	mem(0) := To_stdlogicvector(X"12");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"0A");
	mem(3) := To_stdlogicvector(X"48");
	mem(4) := To_stdlogicvector(X"13");
	mem(5) := To_stdlogicvector(X"66");
	mem(6) := To_stdlogicvector(X"C0");
	mem(7) := To_stdlogicvector(X"40");
	mem(8) := To_stdlogicvector(X"FF");
	mem(9) := To_stdlogicvector(X"0F");
	mem(10) := To_stdlogicvector(X"67");
	mem(11) := To_stdlogicvector(X"12");
	mem(12) := To_stdlogicvector(X"66");
	mem(13) := To_stdlogicvector(X"12");
	mem(14) := To_stdlogicvector(X"65");
	mem(15) := To_stdlogicvector(X"12");
	mem(16) := To_stdlogicvector(X"64");
	mem(17) := To_stdlogicvector(X"12");
	mem(18) := To_stdlogicvector(X"63");
	mem(19) := To_stdlogicvector(X"12");
	mem(20) := To_stdlogicvector(X"62");
	mem(21) := To_stdlogicvector(X"12");
	mem(22) := To_stdlogicvector(X"61");
	mem(23) := To_stdlogicvector(X"12");
	mem(24) := To_stdlogicvector(X"12");
	mem(25) := To_stdlogicvector(X"64");
	mem(26) := To_stdlogicvector(X"25");
	mem(27) := To_stdlogicvector(X"1A");
	mem(28) := To_stdlogicvector(X"C0");
	mem(29) := To_stdlogicvector(X"C1");
	mem(30) := To_stdlogicvector(X"12");
	mem(31) := To_stdlogicvector(X"68");
	mem(32) := To_stdlogicvector(X"26");
	mem(33) := To_stdlogicvector(X"1A");
	mem(34) := To_stdlogicvector(X"C0");
	mem(35) := To_stdlogicvector(X"C1");
	mem(36) := To_stdlogicvector(X"01");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"23");
	mem(39) := To_stdlogicvector(X"00");
