	mem(0) := To_stdlogicvector(X"0A");
	mem(1) := To_stdlogicvector(X"2C");
	mem(2) := To_stdlogicvector(X"0B");
	mem(3) := To_stdlogicvector(X"2E");
	mem(4) := To_stdlogicvector(X"0C");
	mem(5) := To_stdlogicvector(X"3C");
	mem(6) := To_stdlogicvector(X"0D");
	mem(7) := To_stdlogicvector(X"3E");
	mem(8) := To_stdlogicvector(X"FF");
	mem(9) := To_stdlogicvector(X"0F");
	mem(10) := To_stdlogicvector(X"0D");
	mem(11) := To_stdlogicvector(X"60");
	mem(12) := To_stdlogicvector(X"AA");
	mem(13) := To_stdlogicvector(X"BB");
