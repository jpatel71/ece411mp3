	mem(0) := To_stdlogicvector(X"08");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"09");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"0A");
	mem(5) := To_stdlogicvector(X"66");
	mem(6) := To_stdlogicvector(X"63");
	mem(7) := To_stdlogicvector(X"D8");
	mem(8) := To_stdlogicvector(X"98");
	mem(9) := To_stdlogicvector(X"DA");
	mem(10) := To_stdlogicvector(X"B8");
	mem(11) := To_stdlogicvector(X"DC");
	mem(12) := To_stdlogicvector(X"F3");
	mem(13) := To_stdlogicvector(X"DE");
	mem(14) := To_stdlogicvector(X"FF");
	mem(15) := To_stdlogicvector(X"0F");
	mem(16) := To_stdlogicvector(X"01");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"FF");
	mem(19) := To_stdlogicvector(X"FF");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"80");
