LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY ECE411;
USE ECE411.LC3B_TYPES.ALL;

ENTITY MEMORY IS
PORT( 
PMADDRESS  : IN     LC3B_WORD;
PMDATAOUT  : IN     LC3B_OWORD;
PMREAD_L  : IN     STD_LOGIC;
PMWRITE_L : IN     STD_LOGIC;
RESET_L  : IN     STD_LOGIC;
PMDATAIN   : OUT    LC3B_OWORD;
PMRESP_H  : OUT    STD_LOGIC
);
END MEMORY ;

ARCHITECTURE UNTITLED OF MEMORY IS
BEGIN
	-------------------------------------------------------------------
	VHDL_MEMORY : PROCESS (RESET_L, PMREAD_L, PMWRITE_L) 
	-------------------------------------------------------------------
	VARIABLE MEM : MEMORY_ARRAY_64K;
	VARIABLE INT_ADDRESS : INTEGER;
	VARIABLE INT_OLD_ADDRESS : INTEGER;
	BEGIN
		INT_ADDRESS := TO_INTEGER(UNSIGNED(PMADDRESS(12 DOWNTO 4)) * 16);
		IF RESET_L = '0' THEN
			PMRESP_H <= '0';
			MYDRAMINIT_64K(MEM);
		ELSE
			IF ((INT_ADDRESS >= 0) AND (INT_ADDRESS <= 4095)) THEN
				IF (PMWRITE_L'EVENT AND (PMWRITE_L'LAST_VALUE = '0') AND (INT_ADDRESS /= INT_OLD_ADDRESS)) THEN
					ASSERT FALSE 
					REPORT "MEMORY WRITE TIMING ERROR"
					SEVERITY NOTE;
				END IF;
				IF (PMREAD_L'EVENT AND (PMREAD_L'LAST_VALUE = '0') AND (INT_ADDRESS /= INT_OLD_ADDRESS)) THEN
					ASSERT FALSE 
					REPORT "MEMORY READ TIMING ERROR"
					SEVERITY NOTE;
				END IF;
				IF (PMREAD_L = '0' AND PMWRITE_L = '1') THEN
					PMDATAIN(7 DOWNTO 0) <= MEM(INT_ADDRESS) AFTER DELAY_MP22_MEM;            
					PMDATAIN(15 DOWNTO 8) <= MEM(INT_ADDRESS + 1) AFTER DELAY_MP22_MEM;
					PMDATAIN(23 DOWNTO 16) <= MEM(INT_ADDRESS + 2) AFTER DELAY_MP22_MEM;
					PMDATAIN(31 DOWNTO 24) <= MEM(INT_ADDRESS + 3) AFTER DELAY_MP22_MEM;
					PMDATAIN(39 DOWNTO 32) <= MEM(INT_ADDRESS + 4) AFTER DELAY_MP22_MEM;            
					PMDATAIN(47 DOWNTO 40) <= MEM(INT_ADDRESS + 5) AFTER DELAY_MP22_MEM;
					PMDATAIN(55 DOWNTO 48) <= MEM(INT_ADDRESS + 6) AFTER DELAY_MP22_MEM;
					PMDATAIN(63 DOWNTO 56) <= MEM(INT_ADDRESS + 7) AFTER DELAY_MP22_MEM;
					PMDATAIN(71 DOWNTO 64) <= MEM(INT_ADDRESS + 8) AFTER DELAY_MP22_MEM;            
					PMDATAIN(79 DOWNTO 72) <= MEM(INT_ADDRESS + 9) AFTER DELAY_MP22_MEM;
					PMDATAIN(87 DOWNTO 80) <= MEM(INT_ADDRESS + 10) AFTER DELAY_MP22_MEM;
					PMDATAIN(95 DOWNTO 88) <= MEM(INT_ADDRESS + 11) AFTER DELAY_MP22_MEM;
					PMDATAIN(103 DOWNTO 96) <= MEM(INT_ADDRESS + 12) AFTER DELAY_MP22_MEM;            
					PMDATAIN(111 DOWNTO 104) <= MEM(INT_ADDRESS + 13) AFTER DELAY_MP22_MEM;
					PMDATAIN(119 DOWNTO 112) <= MEM(INT_ADDRESS + 14) AFTER DELAY_MP22_MEM;
					PMDATAIN(127 DOWNTO 120) <= MEM(INT_ADDRESS + 15) AFTER DELAY_MP22_MEM;
					PMRESP_H <= '1' AFTER DELAY_MP22_MEM, '0' AFTER (DELAY_MP22_MEM + CLOCK_PERIOD);
				ELSIF (PMWRITE_L = '0' AND PMREAD_L = '1') THEN
					MEM(INT_ADDRESS) := PMDATAOUT(7 DOWNTO 0);
					MEM(INT_ADDRESS + 1) := PMDATAOUT(15 DOWNTO 8);
					MEM(INT_ADDRESS + 2) := PMDATAOUT(23 DOWNTO 16);
					MEM(INT_ADDRESS + 3) := PMDATAOUT(31 DOWNTO 24);
					MEM(INT_ADDRESS + 4) := PMDATAOUT(39 DOWNTO 32);
					MEM(INT_ADDRESS + 5) := PMDATAOUT(47 DOWNTO 40);
					MEM(INT_ADDRESS + 6) := PMDATAOUT(55 DOWNTO 48);
					MEM(INT_ADDRESS + 7) := PMDATAOUT(63 DOWNTO 56);
					MEM(INT_ADDRESS + 8) := PMDATAOUT(71 DOWNTO 64);
					MEM(INT_ADDRESS + 9) := PMDATAOUT(79 DOWNTO 72);
					MEM(INT_ADDRESS + 10) := PMDATAOUT(87 DOWNTO 80);
					MEM(INT_ADDRESS + 11) := PMDATAOUT(95 DOWNTO 88);
					MEM(INT_ADDRESS + 12) := PMDATAOUT(103 DOWNTO 96);
					MEM(INT_ADDRESS + 13) := PMDATAOUT(111 DOWNTO 104);
					MEM(INT_ADDRESS + 14) := PMDATAOUT(119 DOWNTO 112);
					MEM(INT_ADDRESS + 15) := PMDATAOUT(127 DOWNTO 120);
					PMRESP_H <= '1' AFTER DELAY_MP22_MEM, '0' AFTER (DELAY_MP22_MEM + CLOCK_PERIOD);
				ELSE
					ASSERT FALSE 
					REPORT "MEMORY WRITE"
					SEVERITY NOTE;
				END IF;	
			ELSE
				ASSERT FALSE
				REPORT "INVALID ADDRESS"
				SEVERITY WARNING;
			END IF;
		END IF;
	END PROCESS VHDL_MEMORY;
END UNTITLED;
