	mem(0) := To_stdlogicvector(X"21");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"0E");
	mem(3) := To_stdlogicvector(X"0E");
	mem(4) := To_stdlogicvector(X"E7");
	mem(5) := To_stdlogicvector(X"1F");
	mem(6) := To_stdlogicvector(X"E6");
	mem(7) := To_stdlogicvector(X"1F");
	mem(8) := To_stdlogicvector(X"E5");
	mem(9) := To_stdlogicvector(X"1F");
	mem(10) := To_stdlogicvector(X"E4");
	mem(11) := To_stdlogicvector(X"1F");
	mem(12) := To_stdlogicvector(X"21");
	mem(13) := To_stdlogicvector(X"14");
	mem(14) := To_stdlogicvector(X"A2");
	mem(15) := To_stdlogicvector(X"1D");
	mem(16) := To_stdlogicvector(X"FE");
	mem(17) := To_stdlogicvector(X"0F");
	mem(18) := To_stdlogicvector(X"27");
	mem(19) := To_stdlogicvector(X"19");
	mem(20) := To_stdlogicvector(X"26");
	mem(21) := To_stdlogicvector(X"19");
	mem(22) := To_stdlogicvector(X"25");
	mem(23) := To_stdlogicvector(X"19");
	mem(24) := To_stdlogicvector(X"24");
	mem(25) := To_stdlogicvector(X"19");
	mem(26) := To_stdlogicvector(X"23");
	mem(27) := To_stdlogicvector(X"19");
	mem(28) := To_stdlogicvector(X"22");
	mem(29) := To_stdlogicvector(X"19");
	mem(30) := To_stdlogicvector(X"21");
	mem(31) := To_stdlogicvector(X"19");
	mem(32) := To_stdlogicvector(X"25");
	mem(33) := To_stdlogicvector(X"1A");
	mem(34) := To_stdlogicvector(X"F4");
	mem(35) := To_stdlogicvector(X"0F");
