	mem(0) := To_stdlogicvector(X"04");
	mem(1) := To_stdlogicvector(X"AE");
	mem(2) := To_stdlogicvector(X"06");
	mem(3) := To_stdlogicvector(X"BE");
	mem(4) := To_stdlogicvector(X"05");
	mem(5) := To_stdlogicvector(X"68");
	mem(6) := To_stdlogicvector(X"FF");
	mem(7) := To_stdlogicvector(X"0F");
	mem(8) := To_stdlogicvector(X"0A");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"0D");
	mem(11) := To_stdlogicvector(X"60");
	mem(12) := To_stdlogicvector(X"0E");
	mem(13) := To_stdlogicvector(X"00");
