--
-- VHDL Architecture ece411.One.untitled
--
-- Created:
--          by - bjohns38.stdt (eelnx26.ews.illinois.edu)
--          at - 13:41:59 11/10/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.NUMERIC_STD.all;
USE ieee.std_logic_1164.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY One IS
   PORT( 
      clk : IN     std_logic;
      B   : OUT    STD_LOGIC
   );

-- Declarations

END One ;

--
ARCHITECTURE untitled OF One IS
BEGIN
  One<='1';
END ARCHITECTURE untitled;

