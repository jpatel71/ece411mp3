--
-- VHDL Architecture ece411.Adder1.untitled
--
-- Created:
--          by - bjohns38.stdt (eelnx36.ews.illinois.edu)
--          at - 12:28:12 10/18/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.NUMERIC_STD.all;
USE ieee.std_logic_1164.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Adder1 IS
-- Declarations

END Adder1 ;

--
ARCHITECTURE untitled OF Adder1 IS
BEGIN
END ARCHITECTURE untitled;

