ARCHITECTURE UNTITLED OF WORDMUX2 IS
BEGIN
	PROCESS (A, B, SEL)
	VARIABLE STATE : LC3B_WORD;
	BEGIN
		CASE SEL IS
			WHEN '0' =>
				STATE := A;
			WHEN '1' =>
				STATE := B;
			WHEN OTHERS =>
				STATE := (OTHERS => 'X');
		END CASE;
	F <= STATE AFTER DELAY_MUX2;
	END PROCESS;
END UNTITLED;
