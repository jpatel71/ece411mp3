--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - tmurray5.stdt (eelnx33.ews.illinois.edu)
--          at - 15:17:49 08/29/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      ADDRESS   : IN     LC3b_word;
      Clk       : IN     std_logic;
      DATAOUT   : IN     LC3b_word;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      RESET_L   : IN     std_logic;
      DATAIN    : OUT    lc3b_word;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - tmurray5.stdt (eelnx37.ews.illinois.edu)
--          at - 15:42:49 10/14/10
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY ece411;

ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL PMADDRESS    : LC3B_WORD;
   SIGNAL PMDATAIN     : lc3b_oword;
   SIGNAL PMDATAOUT    : LC3B_OWORD;
   SIGNAL PMREAD_L     : STD_LOGIC;
   SIGNAL PMRESP_H     : STD_LOGIC;
   SIGNAL PMWRITE_L    : STD_LOGIC;
   SIGNAL dirty        : std_logic;
   SIGNAL hit          : std_logic;
   SIGNAL in_idleHit   : std_logic;
   SIGNAL in_load      : std_logic;
   SIGNAL in_writeBack : std_logic;
   SIGNAL miss         : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      Clk          : IN     std_logic ;
      PMRESP_H     : IN     STD_LOGIC ;
      RESET_L      : IN     std_logic ;
      dirty        : IN     std_logic ;
      hit          : IN     std_logic ;
      miss         : IN     std_logic ;
      PMREAD_L     : OUT    STD_LOGIC ;
      PMWRITE_L    : OUT    STD_LOGIC ;
      in_idleHit   : OUT    std_logic ;
      in_load      : OUT    std_logic ;
      in_writeBack : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      ADDRESS      : IN     LC3b_word ;
      Clk          : IN     std_logic ;
      DATAOUT      : IN     LC3b_word ;
      MREAD_L      : IN     std_logic ;
      MWRITEH_L    : IN     std_logic ;
      MWRITEL_L    : IN     std_logic ;
      PMDATAIN     : IN     lc3b_oword ;
      RESET_L      : IN     std_logic ;
      in_idleHit   : IN     std_logic ;
      in_load      : IN     std_logic ;
      in_writeback : IN     std_logic ;
      DATAIN       : OUT    lc3b_word ;
      MRESP_H      : OUT    std_logic ;
      PMADDRESS    : OUT    LC3B_WORD ;
      PMDATAOUT    : OUT    lc3b_oword ;
      dirty        : OUT    std_logic ;
      hit          : OUT    std_logic ;
      miss         : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      PMADDRESS : IN     LC3B_WORD ;
      PMREAD_L  : IN     STD_LOGIC ;
      PMWRITE_L : IN     STD_LOGIC ;
      RESET_L   : IN     std_logic ;
      PMDATAIN  : OUT    lc3b_oword ;
      PMRESP_H  : OUT    STD_LOGIC ;
      Clk       : IN     std_logic ;
      PMDATAOUT : IN     LC3B_OWORD 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         Clk          => Clk,
         PMRESP_H     => PMRESP_H,
         RESET_L      => RESET_L,
         dirty        => dirty,
         hit          => hit,
         miss         => miss,
         PMREAD_L     => PMREAD_L,
         PMWRITE_L    => PMWRITE_L,
         in_idleHit   => in_idleHit,
         in_load      => in_load,
         in_writeBack => in_writeBack
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         ADDRESS      => ADDRESS,
         Clk          => Clk,
         DATAOUT      => DATAOUT,
         MREAD_L      => MREAD_L,
         MWRITEH_L    => MWRITEH_L,
         MWRITEL_L    => MWRITEL_L,
         PMDATAIN     => PMDATAIN,
         RESET_L      => RESET_L,
         in_idleHit   => in_idleHit,
         in_load      => in_load,
         in_writeBack => in_writeBack,
         DATAIN       => DATAIN,
         MRESP_H      => MRESP_H,
         PMADDRESS    => PMADDRESS,
         PMDATAOUT    => PMDATAOUT,
         dirty        => dirty,
         hit          => hit,
         miss         => miss
      );
   PDRAM : Physical_Memory
      PORT MAP (
         PMADDRESS => PMADDRESS,
         PMREAD_L  => PMREAD_L,
         PMWRITE_L => PMWRITE_L,
         RESET_L   => RESET_L,
         PMDATAIN  => PMDATAIN,
         PMRESP_H  => PMRESP_H,
         Clk       => Clk,
         PMDATAOUT => PMDATAOUT
      );

END struct;
