	mem(0) := To_stdlogicvector(X"01");
	mem(1) := To_stdlogicvector(X"E2");
	mem(2) := To_stdlogicvector(X"7F");
	mem(3) := To_stdlogicvector(X"94");
	mem(4) := To_stdlogicvector(X"FF");
	mem(5) := To_stdlogicvector(X"0F");
